module top_module( input in, output out );
wire connect;
  assign connect = in;
  assign out = connect;
endmodule
